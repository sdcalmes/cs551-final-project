module cla4(sum, cout, a, b, cin);

input [3:0] a, b;
output [3:0] sum;

input cin;
output cout;

wire [3:0] g, p, c;

//Generate
assign g = a & b;

//Propagate
assign p = a ^ b;

//Carry
assign c[0] = cin;
assign c[1] = g[0] | (p[0] & c[0]);
assign c[2] = g[1] | (p[1] & c[1]);
assign c[3] = g[2] | (p[2] & c[2]);
assign cout = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]) | (p[3] & p[2] & p[1] & p[0] & c[0]);

assign sum = p ^ c;



endmodule

module forwarding(id_rs, id_rt, em_rd, mw_rd, forw_em, forw_mw)
    input [3:0] id_rs, id_rt, em_rd, mw_rd;

endmodule
